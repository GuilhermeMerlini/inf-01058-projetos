library verilog;
use verilog.vl_types.all;
entity Projeto is
    port(
        carga_REM       : out    vl_logic;
        HLT             : out    vl_logic;
        carga_RI        : out    vl_logic;
        clk             : in     vl_logic;
        res             : in     vl_logic;
        RDM_out         : out    vl_logic_vector(7 downto 0);
        read            : out    vl_logic;
        sel             : out    vl_logic;
        PC_out          : out    vl_logic_vector(7 downto 0);
        carga_PC        : out    vl_logic;
        incrementa_PC   : out    vl_logic;
        goto_t0         : out    vl_logic;
        N               : out    vl_logic;
        AC              : out    vl_logic_vector(7 downto 0);
        carga_AC        : out    vl_logic;
        ULA_out         : out    vl_logic_vector(7 downto 0);
        ULAADD          : out    vl_logic;
        ULAAND          : out    vl_logic;
        ULAOR           : out    vl_logic;
        ULANOT          : out    vl_logic;
        ULAy            : out    vl_logic;
        carga_NZ        : out    vl_logic;
        Z               : out    vl_logic;
        NOP             : out    vl_logic;
        STA             : out    vl_logic;
        LDA             : out    vl_logic;
        ADD             : out    vl_logic;
        \OR\            : out    vl_logic;
        \AND\           : out    vl_logic;
        \NOT\           : out    vl_logic;
        JMP             : out    vl_logic;
        JN              : out    vl_logic;
        JZ              : out    vl_logic;
        carga_RDM       : out    vl_logic;
        write           : out    vl_logic;
        ACdisplay0      : out    vl_logic_vector(6 downto 0);
        ACdisplay1      : out    vl_logic_vector(6 downto 0);
        PCdisplay0      : out    vl_logic_vector(6 downto 0);
        PCdisplay1      : out    vl_logic_vector(6 downto 0);
        ROM_out         : out    vl_logic_vector(7 downto 0);
        clk_in          : in     vl_logic
    );
end Projeto;
